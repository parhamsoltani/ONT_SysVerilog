class C4;

endclass