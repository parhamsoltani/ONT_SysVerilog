package param_pkg;

    // global params & typedefs 
    typedef int dimensions_t[2];


    // C4 params & typedefs    
    parameter c4_Length = 260,
              c4_Width = 9, 
              Byte_Num = 8;

    // VC4 params & typedefs
    parameter vc4_Lenght = 261,
              vc4_Width = 9;

    // STM1 params & typedefs          
    parameter STM1_Lenght = 270,
              STM1_Width = 9;


    // CSV params & typedefs
    parameter row_based = 0,
              col_based = 0;


endpackage
