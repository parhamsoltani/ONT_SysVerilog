package class_pkg;
    `include "C4.sv"
endpackage