import param_pkg::*;
import VC4::*;

class AU4;
    VC4 vc4
    byte H1, Y, H2, H3;
    function new();
        vc4 = new();
    endfunction

endclass