package class_pkg;
    `include "C4.sv"
    `include "VC4.sv"
    `include "AU4.sv"
    `include "CSV.sv"
endpackage
