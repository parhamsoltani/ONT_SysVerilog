package param_pkg;

    // global params & typedefs 
    typedef int dimensions_t[2];


    // C4 params & typedefs    
    parameter c4_Length = 260,
              c4_Width = 9, 
              Byte_Num = 8;

    // VC4 params & typedefs    
    parameter vc4_Length = 260,
              vc4_Width = 9;

    // CSV params & typedefs
    parameter row_based = 0,
              col_based = 1;



endpackage