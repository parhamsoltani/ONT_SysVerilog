package class_pkg;
    `include "..\\classes\\C4.sv"
    `include "..\\classes\\VC4.sv"
    `include "..\\classes\\AU4.sv"
    `include "..\\classes\\CSV.sv"
    `include "..\\classes\\STM1.sv"
endpackage
    
