package param_pkg;
    parameter c4_Lenght = 260, c4_Width = 9, Byte_Num = 8 ;
    typedef int c4_index_fixed_array2_t[2];

endpackage