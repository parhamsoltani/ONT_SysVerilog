package param_pkg;

endpackage