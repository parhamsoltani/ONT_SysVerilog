package param_pkg;

    // global params & typedefs 



    // C4 params & typedefs    
    parameter c4_Lenght = 260,
              c4_Width = 9, 
              Byte_Num = 8;

    typedef int c4_index_fixed_array2_t[2];



    // CSV params & typedefs
    parameter row_based = 0,
              col_based = 0;

    typedef int dimensions_t[2];


endpackage
