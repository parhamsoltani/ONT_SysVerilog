package param_pkg;
    parameter c4_Lenght = 260, c4_Width = 9, Byte_Num = 8 ;
    parameter vc4_Lenght = 261, vc4_Width = 9;
    parameter STM1_Lenght = 270, STM1_Width = 9;
    typedef int c4_index_fixed_array2_t[2];

endpackage