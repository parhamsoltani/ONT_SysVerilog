package class_pkg;
    `include "C4.sv"
    `include "VC4.sv"
endpackage