package param_pkg;
    parameter c4_Lenght = 260, c4_Width = 9, Byte_Num = 8 ;
    
    parameter vc4_Lenght = 261, vc4_Width = 9;
    parameter STM1_Lenght = 270, STM1_Width = 9;
    parameter P_letter = 8'b01010000, A_letter = 8'b01000000, R_letter = 8'b01010010, M_letter = 8'b01001101, N_letter = 8'b01001110, SPACE_letter = 8'b00100000;
    typedef int c4_index_fixed_array2_t[2];

endpackage
